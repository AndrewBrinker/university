`include "mod3counter"
`include "adders"
`include "Registers"
`include "instruction_queue"

module tomasulo();


endmodule
