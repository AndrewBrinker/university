module mips();
    // Do the things.
endmodule