`include "test/incr_test.v"
`include "test/mux_test.v"

module test();
    incrTest i();
    muxTest  m();
endmodule
