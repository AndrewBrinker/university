`include "incr_test.v"
`include "mux_test.v"

module test();
    incrTest i();
    muxTest  m();
endmodule
