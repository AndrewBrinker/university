`include "src/fetch/i_fetch.v"
`include "src/decode/i_decode.v"

module pipeline ();



endmodule